

  module inst_mem(CLK, addr, Data,RST);

  input CLK,RST;
  input [5:0]addr;
  output reg[31:0]Data;
  

   always @(*) begin
             case(addr)
	  //******************* reg-reg Operation********************/ 

		 6'd1:    Data =    32'b1100_0100_000011_000100_000101_000000;                 // SUB
                 6'd0:    Data =    32'b1100_0000_000000_000001_000010_000000;                 // ADD               
		 6'd2:    Data =    32'b1100_1000_000110_000111_001000_000000;                 // PASS THROUGH
                 6'd3:    Data =    32'b1100_1100_001001_001010_001011_000000;                 // PASS THROUGH 
		 6'd4:    Data =    32'b1100_0001_001100_001101_001110_000000;                 // LOGICAL AND
	     	 6'd5:    Data =    32'b1100_0101_001111_010000_010001_000000;                 // LOGICAL OR
	         6'd6:    Data =    32'b1100_1001_010010_010011_010100_000000;                 // LOGICAL NOT
		 6'd7:    Data =    32'b1100_1101_010101_010110_010111_000000;                 // LOGICAL EQUALITY
                 6'd8:    Data =    32'b1100_0010_011000_011001_011010_000000;                 // BITWISE AND
		 6'd9:    Data =    32'b1100_0110_011011_011100_011101_000000;                 // BITWISE OR
	        6'd10:    Data =    32'b1100_1010_011110_011111_100000_000000;                 // BITWISE NOT
                6'd11:    Data =    32'b1100_1110_100001_100010_100011_000000;                 // BITWISE XOR             
		6'd12:    Data =    32'b1100_0011_100100_100101_100110_000000;                 // SHIFT RIGHT
	        6'd13:    Data =    32'b1100_0111_100111_101000_101001_000000;                 // SHIFT LEFT
                6'd14:    Data =    32'b1100_1011_101010_101011_101100_000000;                 // ARITHMETIC SHIFT LEFT
                6'd15:    Data =    32'b1100_1111_101101_101110_101111_000000;                 // ARITHMETIC SHIFT RIGHT
		
    
      //********************Reg-Imm Operation********************/ 
 
       6'd17:Data =  32'b1001_0100_000001_000011_1001101011_01;   //SUBI  R3 <- Aimm + R1
       6'd16:Data =  32'b1001_0000_000000_000010_1010100110_01;   // ADDI R2 <- Aimm + R0

      //*****************Imm-reg Instruction*********************/
       
       6'd18: Data = 32'b1010_1001_110100_110101_1011001100_01;  //ORI 
       6'd19: Data = 32'b1110_1000_000110_000111_1010010011_01;  //ANI R7 <- R6 & AIMM
       6'd20: Data = 32'b1101_0010_000000_001011_1010011000_01;  //mov R11 <- AIMM

      //**********************Imm-Imm Instruction***********************//
      
      6'd21:  Data = 32'b1111_0000_101000_01010110_10110010_01; // ADD AIMM Bimm

     //**************************Memory instruction********************************/
      
 
       // Opcode, R_INST, W_INST, ADDR(8(BSEL,REG_SEL+opcode(R_W,X,Y,IN))+ 6 + 6+ 10bit(ADDR) + if(2 bit LSB == 2'b11 then Memory Operation)
       
       // 4 byte
       6'd22: Data = 32'b11_00_1_10_0_000000_001000_0000001100_11; //load  R8 <- data(AX-10)[BSEL+ REG-SEL+ R_W+ X+ Y+ IN+ R_INST+ W_INST+ ADDR+ Memory operation] 
              // 3 byte
       6'd23: Data = 32'b10_00_1_10_0_000000_001100_0000001110_11; //load 
              // 2 byte
       6'd24: Data = 32'b01_00_1_10_0_000000_001001_0000001101_11; //load  
              // 1 byte
       6'd25: Data = 32'b00_00_1_10_0_000000_001001_0000001111_11; //load  
    
       
       //4 byte
       6'd26: Data = 32'b11_00_0_10_0_000100_000000_0010001010_11; //store 
      
       6'd27: Data = 32'b10_00_0_10_0_010100_000000_0011001010_11; //store 
            
       6'd28: Data = 32'b01_00_0_10_0_000110_000000_1010001010_11; //store   
             
       6'd29: Data = 32'b00_00_0_10_0_010101_000000_0010001110_11; //store 
       6'd30: Data = 32'b1101_1100_000000_001011_0000000011_01;    // pass through 
      
       //*******Indirect Addressing Mode******/
        //  CLK --> 1:  Load = R_W=1 + X/Y + IN=1 + R_INST + W_INST
        //  CLK --> 2:  IN=0, R_W=0;
           6'd32: Data = 32'b11_00_1_10_1_001011_011100_0000000000_11;                      
           6'd33: Data = 32'b11_00_0_10_0_001011_011100_0000000000_11;   //Load Operation   

           6'd34: Data = 32'b1101_1100_000000_001111_0000000111_01;      // pass through
	 // Store: CLK --> 1: IN=0, R_INST, R_W=0, X/Y, W_INST(any not required for operation) 
	 //        CLK --> 2: IN=1, R_INST, R_W=0, X/Y, W_INST(any)
        6'd36: Data = 32'b11_00_0_10_0_001111_000000_0000000000_11; 
	6'd37: Data = 32'b11_00_0_10_1_001110_000000_0000000000_11; 
        6'd38: Data = 32'b11_00_1_10_0_000000_000000_0000000001_11;       
      //*********************** Jump Instruction *****************//   
      // {BSEL+REGSEL} + {{X/Y} + R_W + IN} +  ADDR 6 bits + {CON 1 bits + CARRY + PARITY + ZERO} + 2 bits jump op
      //
      //  
      //  Cases:  Absolute jump 
      //          Absolute Conditional Jump
      //          Indirect Jump
      //          Indirect Conditional jump
       
       6'd39:  Data = 32'b1100_010101_010110_010111_000000; 

      6'd40:  Data = 32'b1111_0000_101011_000000000000_0000_10  ; 

       6'd41:  Data = 32'b1111_0000_101100_000000000000_1100_10  ;  // Absolute CON - Carry  
       6'd42:  Data = 32'b1111_0000_101001_000000000000_1010_10  ;  
      6'd43:  Data = 32'b1111_0000_101010_000000000000_1001_10  ; 

      6'd44:  Data = 32'b1111_1011_000010_000000000000_1011_10  ; // Indirect Jump

      6'd46:  Data = 32'b1111_0001_000011_000000000000_1100_10  ; // Indirect CON
      6'd47:  Data = 32'b1111_0001_000100_000000000000_1010_10  ; // Indirect CON
      6'd48:  Data = 32'b1111_0001_000101_000000000000_1001_10  ; // Indirect CON
       

       //*******************  AVERAGE OF 8 NUMBERS *************************//
       // ADD R6,<-- R1, R0
       // ADD R7,<-- R3, R2
       // ADD R8,<-- R5, R4
       // ADD R9,<-- R7, R6
       // ADD R10,<- R6, R7
       // ADD R11,<- R8, R9
       // ADD R12,<- R10, R11
       // Shift_Right A12, Bimm(02)shift right by 2   
      

     /*  6'd49:    Data =    32'b1100_0000_000000_000001_000110_000000;
         6'd50:    Data =    32'b1100_0000_000010_000011_000111_000000;     
         6'd51:    Data =    32'b1100_0000_000100_000101_001000_000000;     
         6'd52:    Data =    32'b1100_0000_000110_000111_001001_000000;     
         6'd53:    Data =    32'b1100_0000_000111_000110_001010_000000;     
         6'd54:    Data =    32'b1100_0000_001001_001000_001011_000000;
         6'd55:    Data =    32'b1100_0000_001011_001010_001100_000000;    */


         6'd49:  Data = 32'b1111_0000_000001_00000010_00000110_01;
         6'd50:  Data = 32'b1111_0000_000010_00000110_00000011_01; 
	 6'd51:  Data = 32'b1111_0000_000011_00000110_00001010_01; 
	 6'd52:  Data = 32'b1111_0000_000100_00001010_00001101_01;

	 6'd53:  Data = 32'b1100_0000_000001_000010_000101_000000;
 	 6'd54:  Data = 32'b1100_0000_000011_000100_000110_000000;

  	 6'd56:  Data = 32'b1100_0000_000110_000101_000111_000000; // add

	 6'd58:  Data =  32'b1101_0011_000111_001000_0000000011_01; // shift

         6'd60:  Data =  32'b1101_0000_001000_001001_0000000000_01; 
	

	  
       
         
	endcase
        end   

	   
	   

	   
endmodule
